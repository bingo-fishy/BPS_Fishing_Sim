module dock_rom
	(
		input wire clk,
		input wire [5:0] row,
		input wire [9:0] col,
		output reg [11:0] color_data
	);

	(* rom_style = "block" *)

	//signal declaration
	reg [5:0] row_reg;
	reg [9:0] col_reg;

	always @(posedge clk)
		begin
		row_reg <= row;
		col_reg <= col;
		end

	always @(*) begin





		if(({row_reg, col_reg}>=16'b0000000000000000) && ({row_reg, col_reg}<16'b0001010000000000)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}>=16'b0001010000000000) && ({row_reg, col_reg}<16'b0001010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001010101100011) && ({row_reg, col_reg}<16'b0001011000111101)) color_data = 12'b000011110000;

		if(({row_reg, col_reg}>=16'b0001011000111101) && ({row_reg, col_reg}<16'b0001100000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100000000000) && ({row_reg, col_reg}<16'b0001100101100011)) color_data = 12'b110110100111;
		if(({row_reg, col_reg}==16'b0001100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001100101100100) && ({row_reg, col_reg}<16'b0001101000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0001101000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0001101000111101) && ({row_reg, col_reg}<16'b0001110101100011)) color_data = 12'b110110100111;
		if(({row_reg, col_reg}==16'b0001110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0001110101100100) && ({row_reg, col_reg}<16'b0001111000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0001111000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0001111000111101) && ({row_reg, col_reg}<16'b0010000101100011)) color_data = 12'b110110100111;
		if(({row_reg, col_reg}==16'b0010000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010000101100100) && ({row_reg, col_reg}<16'b0010001000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0010001000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0010001000111101) && ({row_reg, col_reg}<16'b0010010000000000)) color_data = 12'b110110100111;
		if(({row_reg, col_reg}>=16'b0010010000000000) && ({row_reg, col_reg}<16'b0010010101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0010010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010010101100100) && ({row_reg, col_reg}<16'b0010011000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0010011000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0010011000111101) && ({row_reg, col_reg}<16'b0010100101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0010100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010100101100100) && ({row_reg, col_reg}<16'b0010101000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0010101000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0010101000111101) && ({row_reg, col_reg}<16'b0010110101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0010110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0010110101100100) && ({row_reg, col_reg}<16'b0010111000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0010111000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0010111000111101) && ({row_reg, col_reg}<16'b0011000101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0011000101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011000101100100) && ({row_reg, col_reg}<16'b0011001000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0011001000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011001000111101) && ({row_reg, col_reg}<16'b0011010101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0011010101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011010101100100) && ({row_reg, col_reg}<16'b0011011000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0011011000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011011000111101) && ({row_reg, col_reg}<16'b0011100101100011)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}==16'b0011100101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011100101100100) && ({row_reg, col_reg}<16'b0011101000111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0011101000111100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0011101000111101) && ({row_reg, col_reg}<16'b0011110000000000)) color_data = 12'b110110010101;
		if(({row_reg, col_reg}>=16'b0011110000000000) && ({row_reg, col_reg}<16'b0011110000011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110000011010) && ({row_reg, col_reg}<16'b0011110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0011110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}>=16'b0011110000101010) && ({row_reg, col_reg}<16'b0011110001111110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110001111110) && ({row_reg, col_reg}<16'b0011110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0011110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}>=16'b0011110010001110) && ({row_reg, col_reg}<16'b0011110011011110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110011011110) && ({row_reg, col_reg}<16'b0011110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}>=16'b0011110011101101) && ({row_reg, col_reg}<16'b0011110101000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110101000000) && ({row_reg, col_reg}<16'b0011110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}>=16'b0011110101001111) && ({row_reg, col_reg}<16'b0011110101100011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011110101100011) && ({row_reg, col_reg}<16'b0011111000111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}>=16'b0011111000111101) && ({row_reg, col_reg}<16'b0011111001010111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111001010111) && ({row_reg, col_reg}<16'b0011111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0011111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}>=16'b0011111001100111) && ({row_reg, col_reg}<16'b0011111010111011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111010111011) && ({row_reg, col_reg}<16'b0011111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0011111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}>=16'b0011111011001011) && ({row_reg, col_reg}<16'b0011111100011011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111100011011) && ({row_reg, col_reg}<16'b0011111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}>=16'b0011111100101010) && ({row_reg, col_reg}<16'b0011111101111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0011111101111101) && ({row_reg, col_reg}<16'b0011111110001100)) color_data = 12'b101101110011;

		if(({row_reg, col_reg}>=16'b0011111110001100) && ({row_reg, col_reg}<16'b0100000000000000)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000000000) && ({row_reg, col_reg}<16'b0100000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000011010) && ({row_reg, col_reg}<16'b0100000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000000101011) && ({row_reg, col_reg}<16'b0100000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000001111110) && ({row_reg, col_reg}<16'b0100000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000010001111) && ({row_reg, col_reg}<16'b0100000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000011011110) && ({row_reg, col_reg}<16'b0100000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000011101110) && ({row_reg, col_reg}<16'b0100000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000101000000) && ({row_reg, col_reg}<16'b0100000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100000101010000) && ({row_reg, col_reg}<16'b0100001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001001010111) && ({row_reg, col_reg}<16'b0100001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001001101000) && ({row_reg, col_reg}<16'b0100001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001010111011) && ({row_reg, col_reg}<16'b0100001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001011001100) && ({row_reg, col_reg}<16'b0100001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100011011) && ({row_reg, col_reg}<16'b0100001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001100101011) && ({row_reg, col_reg}<16'b0100001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100001101111101) && ({row_reg, col_reg}<16'b0100001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100001110001101) && ({row_reg, col_reg}<16'b0100010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010000011010) && ({row_reg, col_reg}<16'b0100010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010000101011) && ({row_reg, col_reg}<16'b0100010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010001111110) && ({row_reg, col_reg}<16'b0100010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010010001111) && ({row_reg, col_reg}<16'b0100010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010011011110) && ({row_reg, col_reg}<16'b0100010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010011101110) && ({row_reg, col_reg}<16'b0100010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010101000000) && ({row_reg, col_reg}<16'b0100010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100010101010000) && ({row_reg, col_reg}<16'b0100011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011001010111) && ({row_reg, col_reg}<16'b0100011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011001101000) && ({row_reg, col_reg}<16'b0100011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011010111011) && ({row_reg, col_reg}<16'b0100011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011011001100) && ({row_reg, col_reg}<16'b0100011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011100011011) && ({row_reg, col_reg}<16'b0100011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011100101011) && ({row_reg, col_reg}<16'b0100011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100011101111101) && ({row_reg, col_reg}<16'b0100011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100011110001101) && ({row_reg, col_reg}<16'b0100100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100000011010) && ({row_reg, col_reg}<16'b0100100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100000101011) && ({row_reg, col_reg}<16'b0100100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100001111110) && ({row_reg, col_reg}<16'b0100100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100010001111) && ({row_reg, col_reg}<16'b0100100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100011011110) && ({row_reg, col_reg}<16'b0100100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100011101110) && ({row_reg, col_reg}<16'b0100100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100101000000) && ({row_reg, col_reg}<16'b0100100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100100101010000) && ({row_reg, col_reg}<16'b0100101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101001010111) && ({row_reg, col_reg}<16'b0100101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101001101000) && ({row_reg, col_reg}<16'b0100101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101010111011) && ({row_reg, col_reg}<16'b0100101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101011001100) && ({row_reg, col_reg}<16'b0100101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101100011011) && ({row_reg, col_reg}<16'b0100101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101100101011) && ({row_reg, col_reg}<16'b0100101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100101101111101) && ({row_reg, col_reg}<16'b0100101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100101110001101) && ({row_reg, col_reg}<16'b0100110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110000011010) && ({row_reg, col_reg}<16'b0100110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110000101011) && ({row_reg, col_reg}<16'b0100110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110001111110) && ({row_reg, col_reg}<16'b0100110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110010001111) && ({row_reg, col_reg}<16'b0100110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110011011110) && ({row_reg, col_reg}<16'b0100110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110011101110) && ({row_reg, col_reg}<16'b0100110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110101000000) && ({row_reg, col_reg}<16'b0100110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100110101010000) && ({row_reg, col_reg}<16'b0100111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111001010111) && ({row_reg, col_reg}<16'b0100111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0100111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111001101000) && ({row_reg, col_reg}<16'b0100111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111010111011) && ({row_reg, col_reg}<16'b0100111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0100111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111011001100) && ({row_reg, col_reg}<16'b0100111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111100011011) && ({row_reg, col_reg}<16'b0100111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111100101011) && ({row_reg, col_reg}<16'b0100111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0100111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0100111101111101) && ({row_reg, col_reg}<16'b0100111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0100111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0100111110001101) && ({row_reg, col_reg}<16'b0101000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000000011010) && ({row_reg, col_reg}<16'b0101000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000000101011) && ({row_reg, col_reg}<16'b0101000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000001111110) && ({row_reg, col_reg}<16'b0101000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000010001111) && ({row_reg, col_reg}<16'b0101000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000011011110) && ({row_reg, col_reg}<16'b0101000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000011101110) && ({row_reg, col_reg}<16'b0101000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000101000000) && ({row_reg, col_reg}<16'b0101000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101000101010000) && ({row_reg, col_reg}<16'b0101001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001001010111) && ({row_reg, col_reg}<16'b0101001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001001101000) && ({row_reg, col_reg}<16'b0101001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001010111011) && ({row_reg, col_reg}<16'b0101001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001011001100) && ({row_reg, col_reg}<16'b0101001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001100011011) && ({row_reg, col_reg}<16'b0101001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001100101011) && ({row_reg, col_reg}<16'b0101001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101001101111101) && ({row_reg, col_reg}<16'b0101001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101001110001101) && ({row_reg, col_reg}<16'b0101010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010000011010) && ({row_reg, col_reg}<16'b0101010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010000101011) && ({row_reg, col_reg}<16'b0101010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010001111110) && ({row_reg, col_reg}<16'b0101010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010010001111) && ({row_reg, col_reg}<16'b0101010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011011110) && ({row_reg, col_reg}<16'b0101010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010011101110) && ({row_reg, col_reg}<16'b0101010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010101000000) && ({row_reg, col_reg}<16'b0101010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101010101010000) && ({row_reg, col_reg}<16'b0101011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011001010111) && ({row_reg, col_reg}<16'b0101011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011001101000) && ({row_reg, col_reg}<16'b0101011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011010111011) && ({row_reg, col_reg}<16'b0101011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011011001100) && ({row_reg, col_reg}<16'b0101011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011100011011) && ({row_reg, col_reg}<16'b0101011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011100101011) && ({row_reg, col_reg}<16'b0101011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101011101111101) && ({row_reg, col_reg}<16'b0101011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101011110001101) && ({row_reg, col_reg}<16'b0101100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100000011010) && ({row_reg, col_reg}<16'b0101100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100000101011) && ({row_reg, col_reg}<16'b0101100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100001111110) && ({row_reg, col_reg}<16'b0101100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100010001111) && ({row_reg, col_reg}<16'b0101100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100011011110) && ({row_reg, col_reg}<16'b0101100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100011101110) && ({row_reg, col_reg}<16'b0101100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100101000000) && ({row_reg, col_reg}<16'b0101100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101100101010000) && ({row_reg, col_reg}<16'b0101101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101001010111) && ({row_reg, col_reg}<16'b0101101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101001101000) && ({row_reg, col_reg}<16'b0101101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101010111011) && ({row_reg, col_reg}<16'b0101101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101011001100) && ({row_reg, col_reg}<16'b0101101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101100011011) && ({row_reg, col_reg}<16'b0101101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101100101011) && ({row_reg, col_reg}<16'b0101101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101101101111101) && ({row_reg, col_reg}<16'b0101101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101101110001101) && ({row_reg, col_reg}<16'b0101110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110000011010) && ({row_reg, col_reg}<16'b0101110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110000101011) && ({row_reg, col_reg}<16'b0101110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110001111110) && ({row_reg, col_reg}<16'b0101110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110010001111) && ({row_reg, col_reg}<16'b0101110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110011011110) && ({row_reg, col_reg}<16'b0101110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110011101110) && ({row_reg, col_reg}<16'b0101110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110101000000) && ({row_reg, col_reg}<16'b0101110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101110101010000) && ({row_reg, col_reg}<16'b0101111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111001010111) && ({row_reg, col_reg}<16'b0101111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0101111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111001101000) && ({row_reg, col_reg}<16'b0101111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111010111011) && ({row_reg, col_reg}<16'b0101111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0101111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111011001100) && ({row_reg, col_reg}<16'b0101111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111100011011) && ({row_reg, col_reg}<16'b0101111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111100101011) && ({row_reg, col_reg}<16'b0101111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0101111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0101111101111101) && ({row_reg, col_reg}<16'b0101111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0101111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0101111110001101) && ({row_reg, col_reg}<16'b0110000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000000011010) && ({row_reg, col_reg}<16'b0110000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000000101011) && ({row_reg, col_reg}<16'b0110000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000001111110) && ({row_reg, col_reg}<16'b0110000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000010001111) && ({row_reg, col_reg}<16'b0110000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000011011110) && ({row_reg, col_reg}<16'b0110000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000011101110) && ({row_reg, col_reg}<16'b0110000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000101000000) && ({row_reg, col_reg}<16'b0110000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110000101010000) && ({row_reg, col_reg}<16'b0110001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001001010111) && ({row_reg, col_reg}<16'b0110001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001001101000) && ({row_reg, col_reg}<16'b0110001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001010111011) && ({row_reg, col_reg}<16'b0110001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001011001100) && ({row_reg, col_reg}<16'b0110001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001100011011) && ({row_reg, col_reg}<16'b0110001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001100101011) && ({row_reg, col_reg}<16'b0110001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110001101111101) && ({row_reg, col_reg}<16'b0110001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0110001110001101) && ({row_reg, col_reg}<16'b0110010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010000011010) && ({row_reg, col_reg}<16'b0110010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010000101011) && ({row_reg, col_reg}<16'b0110010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010001111110) && ({row_reg, col_reg}<16'b0110010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010010001111) && ({row_reg, col_reg}<16'b0110010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011011110) && ({row_reg, col_reg}<16'b0110010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010011101110) && ({row_reg, col_reg}<16'b0110010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010101000000) && ({row_reg, col_reg}<16'b0110010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110010101010000) && ({row_reg, col_reg}<16'b0110011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011001010111) && ({row_reg, col_reg}<16'b0110011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011001101000) && ({row_reg, col_reg}<16'b0110011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011010111011) && ({row_reg, col_reg}<16'b0110011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011011001100) && ({row_reg, col_reg}<16'b0110011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011100011011) && ({row_reg, col_reg}<16'b0110011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011100101011) && ({row_reg, col_reg}<16'b0110011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110011101111101) && ({row_reg, col_reg}<16'b0110011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0110011110001101) && ({row_reg, col_reg}<16'b0110100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100000011010) && ({row_reg, col_reg}<16'b0110100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100000101011) && ({row_reg, col_reg}<16'b0110100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100001111110) && ({row_reg, col_reg}<16'b0110100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100010001111) && ({row_reg, col_reg}<16'b0110100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100011011110) && ({row_reg, col_reg}<16'b0110100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100011101110) && ({row_reg, col_reg}<16'b0110100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100101000000) && ({row_reg, col_reg}<16'b0110100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110100101010000) && ({row_reg, col_reg}<16'b0110101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101001010111) && ({row_reg, col_reg}<16'b0110101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101001101000) && ({row_reg, col_reg}<16'b0110101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101010111011) && ({row_reg, col_reg}<16'b0110101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101011001100) && ({row_reg, col_reg}<16'b0110101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101100011011) && ({row_reg, col_reg}<16'b0110101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101100101011) && ({row_reg, col_reg}<16'b0110101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110101101111101) && ({row_reg, col_reg}<16'b0110101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0110101110001101) && ({row_reg, col_reg}<16'b0110110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110000011010) && ({row_reg, col_reg}<16'b0110110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110000101011) && ({row_reg, col_reg}<16'b0110110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110001111110) && ({row_reg, col_reg}<16'b0110110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110010001111) && ({row_reg, col_reg}<16'b0110110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110011011110) && ({row_reg, col_reg}<16'b0110110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110011101110) && ({row_reg, col_reg}<16'b0110110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110101000000) && ({row_reg, col_reg}<16'b0110110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110110101010000) && ({row_reg, col_reg}<16'b0110111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111001010111) && ({row_reg, col_reg}<16'b0110111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0110111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111001101000) && ({row_reg, col_reg}<16'b0110111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111010111011) && ({row_reg, col_reg}<16'b0110111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0110111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111011001100) && ({row_reg, col_reg}<16'b0110111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111100011011) && ({row_reg, col_reg}<16'b0110111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111100101011) && ({row_reg, col_reg}<16'b0110111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0110111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0110111101111101) && ({row_reg, col_reg}<16'b0110111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0110111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0110111110001101) && ({row_reg, col_reg}<16'b0111000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000011010) && ({row_reg, col_reg}<16'b0111000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000000101011) && ({row_reg, col_reg}<16'b0111000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000001111110) && ({row_reg, col_reg}<16'b0111000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000010001111) && ({row_reg, col_reg}<16'b0111000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000011011110) && ({row_reg, col_reg}<16'b0111000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000011101110) && ({row_reg, col_reg}<16'b0111000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000101000000) && ({row_reg, col_reg}<16'b0111000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111000101010000) && ({row_reg, col_reg}<16'b0111001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001001010111) && ({row_reg, col_reg}<16'b0111001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001001101000) && ({row_reg, col_reg}<16'b0111001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001010111011) && ({row_reg, col_reg}<16'b0111001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001011001100) && ({row_reg, col_reg}<16'b0111001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001100011011) && ({row_reg, col_reg}<16'b0111001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001100101011) && ({row_reg, col_reg}<16'b0111001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111001101111101) && ({row_reg, col_reg}<16'b0111001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111001110001101) && ({row_reg, col_reg}<16'b0111010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010000011010) && ({row_reg, col_reg}<16'b0111010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010000101011) && ({row_reg, col_reg}<16'b0111010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010001111110) && ({row_reg, col_reg}<16'b0111010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010010001111) && ({row_reg, col_reg}<16'b0111010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010011011110) && ({row_reg, col_reg}<16'b0111010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010011101110) && ({row_reg, col_reg}<16'b0111010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010101000000) && ({row_reg, col_reg}<16'b0111010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111010101010000) && ({row_reg, col_reg}<16'b0111011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011001010111) && ({row_reg, col_reg}<16'b0111011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011001101000) && ({row_reg, col_reg}<16'b0111011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011010111011) && ({row_reg, col_reg}<16'b0111011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011011001100) && ({row_reg, col_reg}<16'b0111011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011100011011) && ({row_reg, col_reg}<16'b0111011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011100101011) && ({row_reg, col_reg}<16'b0111011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111011101111101) && ({row_reg, col_reg}<16'b0111011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111011110001101) && ({row_reg, col_reg}<16'b0111100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100000011010) && ({row_reg, col_reg}<16'b0111100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100000101011) && ({row_reg, col_reg}<16'b0111100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100001111110) && ({row_reg, col_reg}<16'b0111100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100010001111) && ({row_reg, col_reg}<16'b0111100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100011011110) && ({row_reg, col_reg}<16'b0111100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100011101110) && ({row_reg, col_reg}<16'b0111100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100101000000) && ({row_reg, col_reg}<16'b0111100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111100101010000) && ({row_reg, col_reg}<16'b0111101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101001010111) && ({row_reg, col_reg}<16'b0111101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101001101000) && ({row_reg, col_reg}<16'b0111101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101010111011) && ({row_reg, col_reg}<16'b0111101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101011001100) && ({row_reg, col_reg}<16'b0111101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101100011011) && ({row_reg, col_reg}<16'b0111101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101100101011) && ({row_reg, col_reg}<16'b0111101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111101101111101) && ({row_reg, col_reg}<16'b0111101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111101110001101) && ({row_reg, col_reg}<16'b0111110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000011010) && ({row_reg, col_reg}<16'b0111110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110000101011) && ({row_reg, col_reg}<16'b0111110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110001111110) && ({row_reg, col_reg}<16'b0111110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110010001111) && ({row_reg, col_reg}<16'b0111110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110011011110) && ({row_reg, col_reg}<16'b0111110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110011101110) && ({row_reg, col_reg}<16'b0111110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110101000000) && ({row_reg, col_reg}<16'b0111110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111110101010000) && ({row_reg, col_reg}<16'b0111111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111001010111) && ({row_reg, col_reg}<16'b0111111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b0111111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111001101000) && ({row_reg, col_reg}<16'b0111111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111010111011) && ({row_reg, col_reg}<16'b0111111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b0111111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111011001100) && ({row_reg, col_reg}<16'b0111111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111100011011) && ({row_reg, col_reg}<16'b0111111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111100101011) && ({row_reg, col_reg}<16'b0111111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b0111111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b0111111101111101) && ({row_reg, col_reg}<16'b0111111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b0111111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b0111111110001101) && ({row_reg, col_reg}<16'b1000000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000000011010) && ({row_reg, col_reg}<16'b1000000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000000101011) && ({row_reg, col_reg}<16'b1000000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000001111110) && ({row_reg, col_reg}<16'b1000000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000010001111) && ({row_reg, col_reg}<16'b1000000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000011011110) && ({row_reg, col_reg}<16'b1000000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000011101110) && ({row_reg, col_reg}<16'b1000000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000101000000) && ({row_reg, col_reg}<16'b1000000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000000101010000) && ({row_reg, col_reg}<16'b1000001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001001010111) && ({row_reg, col_reg}<16'b1000001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001001101000) && ({row_reg, col_reg}<16'b1000001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001010111011) && ({row_reg, col_reg}<16'b1000001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001011001100) && ({row_reg, col_reg}<16'b1000001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001100011011) && ({row_reg, col_reg}<16'b1000001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001100101011) && ({row_reg, col_reg}<16'b1000001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000001101111101) && ({row_reg, col_reg}<16'b1000001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000001110001101) && ({row_reg, col_reg}<16'b1000010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010000011010) && ({row_reg, col_reg}<16'b1000010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010000101011) && ({row_reg, col_reg}<16'b1000010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010001111110) && ({row_reg, col_reg}<16'b1000010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010010001111) && ({row_reg, col_reg}<16'b1000010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010011011110) && ({row_reg, col_reg}<16'b1000010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010011101110) && ({row_reg, col_reg}<16'b1000010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010101000000) && ({row_reg, col_reg}<16'b1000010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000010101010000) && ({row_reg, col_reg}<16'b1000011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011001010111) && ({row_reg, col_reg}<16'b1000011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011001101000) && ({row_reg, col_reg}<16'b1000011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011010111011) && ({row_reg, col_reg}<16'b1000011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011011001100) && ({row_reg, col_reg}<16'b1000011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011100011011) && ({row_reg, col_reg}<16'b1000011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011100101011) && ({row_reg, col_reg}<16'b1000011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000011101111101) && ({row_reg, col_reg}<16'b1000011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000011110001101) && ({row_reg, col_reg}<16'b1000100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100000011010) && ({row_reg, col_reg}<16'b1000100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100000101011) && ({row_reg, col_reg}<16'b1000100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100001111110) && ({row_reg, col_reg}<16'b1000100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100010001111) && ({row_reg, col_reg}<16'b1000100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100011011110) && ({row_reg, col_reg}<16'b1000100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100011101110) && ({row_reg, col_reg}<16'b1000100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100101000000) && ({row_reg, col_reg}<16'b1000100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000100101010000) && ({row_reg, col_reg}<16'b1000101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101001010111) && ({row_reg, col_reg}<16'b1000101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101001101000) && ({row_reg, col_reg}<16'b1000101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101010111011) && ({row_reg, col_reg}<16'b1000101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101011001100) && ({row_reg, col_reg}<16'b1000101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101100011011) && ({row_reg, col_reg}<16'b1000101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101100101011) && ({row_reg, col_reg}<16'b1000101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000101101111101) && ({row_reg, col_reg}<16'b1000101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000101110001101) && ({row_reg, col_reg}<16'b1000110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110000011010) && ({row_reg, col_reg}<16'b1000110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110000101011) && ({row_reg, col_reg}<16'b1000110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110001111110) && ({row_reg, col_reg}<16'b1000110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110010001111) && ({row_reg, col_reg}<16'b1000110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110011011110) && ({row_reg, col_reg}<16'b1000110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110011101110) && ({row_reg, col_reg}<16'b1000110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110101000000) && ({row_reg, col_reg}<16'b1000110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000110101010000) && ({row_reg, col_reg}<16'b1000111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111001010111) && ({row_reg, col_reg}<16'b1000111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1000111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111001101000) && ({row_reg, col_reg}<16'b1000111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111010111011) && ({row_reg, col_reg}<16'b1000111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1000111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111011001100) && ({row_reg, col_reg}<16'b1000111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111100011011) && ({row_reg, col_reg}<16'b1000111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111100101011) && ({row_reg, col_reg}<16'b1000111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1000111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1000111101111101) && ({row_reg, col_reg}<16'b1000111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1000111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1000111110001101) && ({row_reg, col_reg}<16'b1001000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000000011010) && ({row_reg, col_reg}<16'b1001000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000000101011) && ({row_reg, col_reg}<16'b1001000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000001111110) && ({row_reg, col_reg}<16'b1001000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000010001111) && ({row_reg, col_reg}<16'b1001000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000011011110) && ({row_reg, col_reg}<16'b1001000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000011101110) && ({row_reg, col_reg}<16'b1001000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000101000000) && ({row_reg, col_reg}<16'b1001000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001000101010000) && ({row_reg, col_reg}<16'b1001001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001001010111) && ({row_reg, col_reg}<16'b1001001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001001101000) && ({row_reg, col_reg}<16'b1001001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001010111011) && ({row_reg, col_reg}<16'b1001001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001011001100) && ({row_reg, col_reg}<16'b1001001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001100011011) && ({row_reg, col_reg}<16'b1001001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001100101011) && ({row_reg, col_reg}<16'b1001001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001001101111101) && ({row_reg, col_reg}<16'b1001001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1001001110001101) && ({row_reg, col_reg}<16'b1001010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010000011010) && ({row_reg, col_reg}<16'b1001010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010000101011) && ({row_reg, col_reg}<16'b1001010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010001111110) && ({row_reg, col_reg}<16'b1001010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010010001111) && ({row_reg, col_reg}<16'b1001010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010011011110) && ({row_reg, col_reg}<16'b1001010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010011101110) && ({row_reg, col_reg}<16'b1001010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010101000000) && ({row_reg, col_reg}<16'b1001010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001010101010000) && ({row_reg, col_reg}<16'b1001011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011001010111) && ({row_reg, col_reg}<16'b1001011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011001101000) && ({row_reg, col_reg}<16'b1001011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011010111011) && ({row_reg, col_reg}<16'b1001011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011011001100) && ({row_reg, col_reg}<16'b1001011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011100011011) && ({row_reg, col_reg}<16'b1001011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011100101011) && ({row_reg, col_reg}<16'b1001011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001011101111101) && ({row_reg, col_reg}<16'b1001011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1001011110001101) && ({row_reg, col_reg}<16'b1001100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100000011010) && ({row_reg, col_reg}<16'b1001100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100000101011) && ({row_reg, col_reg}<16'b1001100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100001111110) && ({row_reg, col_reg}<16'b1001100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100010001111) && ({row_reg, col_reg}<16'b1001100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100011011110) && ({row_reg, col_reg}<16'b1001100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100011101110) && ({row_reg, col_reg}<16'b1001100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100101000000) && ({row_reg, col_reg}<16'b1001100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001100101010000) && ({row_reg, col_reg}<16'b1001101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101001010111) && ({row_reg, col_reg}<16'b1001101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101001101000) && ({row_reg, col_reg}<16'b1001101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101010111011) && ({row_reg, col_reg}<16'b1001101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101011001100) && ({row_reg, col_reg}<16'b1001101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101100011011) && ({row_reg, col_reg}<16'b1001101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101100101011) && ({row_reg, col_reg}<16'b1001101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001101101111101) && ({row_reg, col_reg}<16'b1001101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1001101110001101) && ({row_reg, col_reg}<16'b1001110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110000011010) && ({row_reg, col_reg}<16'b1001110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110000101011) && ({row_reg, col_reg}<16'b1001110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110001111110) && ({row_reg, col_reg}<16'b1001110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110010001111) && ({row_reg, col_reg}<16'b1001110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110011011110) && ({row_reg, col_reg}<16'b1001110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110011101110) && ({row_reg, col_reg}<16'b1001110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110101000000) && ({row_reg, col_reg}<16'b1001110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001110101010000) && ({row_reg, col_reg}<16'b1001111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111001010111) && ({row_reg, col_reg}<16'b1001111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1001111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111001101000) && ({row_reg, col_reg}<16'b1001111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111010111011) && ({row_reg, col_reg}<16'b1001111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1001111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111011001100) && ({row_reg, col_reg}<16'b1001111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111100011011) && ({row_reg, col_reg}<16'b1001111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111100101011) && ({row_reg, col_reg}<16'b1001111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1001111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1001111101111101) && ({row_reg, col_reg}<16'b1001111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1001111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1001111110001101) && ({row_reg, col_reg}<16'b1010000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000000011010) && ({row_reg, col_reg}<16'b1010000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000000101011) && ({row_reg, col_reg}<16'b1010000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000001111110) && ({row_reg, col_reg}<16'b1010000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000010001111) && ({row_reg, col_reg}<16'b1010000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000011011110) && ({row_reg, col_reg}<16'b1010000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000011101110) && ({row_reg, col_reg}<16'b1010000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000101000000) && ({row_reg, col_reg}<16'b1010000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010000101010000) && ({row_reg, col_reg}<16'b1010001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001001010111) && ({row_reg, col_reg}<16'b1010001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001001101000) && ({row_reg, col_reg}<16'b1010001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001010111011) && ({row_reg, col_reg}<16'b1010001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001011001100) && ({row_reg, col_reg}<16'b1010001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001100011011) && ({row_reg, col_reg}<16'b1010001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001100101011) && ({row_reg, col_reg}<16'b1010001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010001101111101) && ({row_reg, col_reg}<16'b1010001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1010001110001101) && ({row_reg, col_reg}<16'b1010010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010000011010) && ({row_reg, col_reg}<16'b1010010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010000101011) && ({row_reg, col_reg}<16'b1010010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010001111110) && ({row_reg, col_reg}<16'b1010010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010010001111) && ({row_reg, col_reg}<16'b1010010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010011011110) && ({row_reg, col_reg}<16'b1010010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010011101110) && ({row_reg, col_reg}<16'b1010010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010101000000) && ({row_reg, col_reg}<16'b1010010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010010101010000) && ({row_reg, col_reg}<16'b1010011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011001010111) && ({row_reg, col_reg}<16'b1010011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011001101000) && ({row_reg, col_reg}<16'b1010011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011010111011) && ({row_reg, col_reg}<16'b1010011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011011001100) && ({row_reg, col_reg}<16'b1010011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011100011011) && ({row_reg, col_reg}<16'b1010011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011100101011) && ({row_reg, col_reg}<16'b1010011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010011101111101) && ({row_reg, col_reg}<16'b1010011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1010011110001101) && ({row_reg, col_reg}<16'b1010100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100000011010) && ({row_reg, col_reg}<16'b1010100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100000101011) && ({row_reg, col_reg}<16'b1010100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100001111110) && ({row_reg, col_reg}<16'b1010100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100010001111) && ({row_reg, col_reg}<16'b1010100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100011011110) && ({row_reg, col_reg}<16'b1010100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100011101110) && ({row_reg, col_reg}<16'b1010100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100101000000) && ({row_reg, col_reg}<16'b1010100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010100101010000) && ({row_reg, col_reg}<16'b1010101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101001010111) && ({row_reg, col_reg}<16'b1010101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101001101000) && ({row_reg, col_reg}<16'b1010101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101010111011) && ({row_reg, col_reg}<16'b1010101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101011001100) && ({row_reg, col_reg}<16'b1010101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101100011011) && ({row_reg, col_reg}<16'b1010101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101100101011) && ({row_reg, col_reg}<16'b1010101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010101101111101) && ({row_reg, col_reg}<16'b1010101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1010101110001101) && ({row_reg, col_reg}<16'b1010110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110000011010) && ({row_reg, col_reg}<16'b1010110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110000101011) && ({row_reg, col_reg}<16'b1010110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110001111110) && ({row_reg, col_reg}<16'b1010110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110010001111) && ({row_reg, col_reg}<16'b1010110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110011011110) && ({row_reg, col_reg}<16'b1010110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110011101110) && ({row_reg, col_reg}<16'b1010110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110101000000) && ({row_reg, col_reg}<16'b1010110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010110101010000) && ({row_reg, col_reg}<16'b1010111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111001010111) && ({row_reg, col_reg}<16'b1010111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1010111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111001101000) && ({row_reg, col_reg}<16'b1010111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111010111011) && ({row_reg, col_reg}<16'b1010111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1010111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111011001100) && ({row_reg, col_reg}<16'b1010111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111100011011) && ({row_reg, col_reg}<16'b1010111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111100101011) && ({row_reg, col_reg}<16'b1010111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1010111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1010111101111101) && ({row_reg, col_reg}<16'b1010111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1010111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1010111110001101) && ({row_reg, col_reg}<16'b1011000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000000011010) && ({row_reg, col_reg}<16'b1011000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000000101011) && ({row_reg, col_reg}<16'b1011000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000001111110) && ({row_reg, col_reg}<16'b1011000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000010001111) && ({row_reg, col_reg}<16'b1011000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000011011110) && ({row_reg, col_reg}<16'b1011000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000011101110) && ({row_reg, col_reg}<16'b1011000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000101000000) && ({row_reg, col_reg}<16'b1011000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011000101010000) && ({row_reg, col_reg}<16'b1011001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001001010111) && ({row_reg, col_reg}<16'b1011001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001001101000) && ({row_reg, col_reg}<16'b1011001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001010111011) && ({row_reg, col_reg}<16'b1011001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001011001100) && ({row_reg, col_reg}<16'b1011001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001100011011) && ({row_reg, col_reg}<16'b1011001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001100101011) && ({row_reg, col_reg}<16'b1011001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011001101111101) && ({row_reg, col_reg}<16'b1011001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1011001110001101) && ({row_reg, col_reg}<16'b1011010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010000011010) && ({row_reg, col_reg}<16'b1011010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010000101011) && ({row_reg, col_reg}<16'b1011010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010001111110) && ({row_reg, col_reg}<16'b1011010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010010001111) && ({row_reg, col_reg}<16'b1011010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010011011110) && ({row_reg, col_reg}<16'b1011010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010011101110) && ({row_reg, col_reg}<16'b1011010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010101000000) && ({row_reg, col_reg}<16'b1011010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011010101010000) && ({row_reg, col_reg}<16'b1011011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011001010111) && ({row_reg, col_reg}<16'b1011011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011001101000) && ({row_reg, col_reg}<16'b1011011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011010111011) && ({row_reg, col_reg}<16'b1011011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011011001100) && ({row_reg, col_reg}<16'b1011011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011100011011) && ({row_reg, col_reg}<16'b1011011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011100101011) && ({row_reg, col_reg}<16'b1011011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011011101111101) && ({row_reg, col_reg}<16'b1011011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1011011110001101) && ({row_reg, col_reg}<16'b1011100000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011100000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100000011010) && ({row_reg, col_reg}<16'b1011100000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011100000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011100000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100000101011) && ({row_reg, col_reg}<16'b1011100001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011100001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100001111110) && ({row_reg, col_reg}<16'b1011100010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011100010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011100010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100010001111) && ({row_reg, col_reg}<16'b1011100011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011100011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100011011110) && ({row_reg, col_reg}<16'b1011100011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011100011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100011101110) && ({row_reg, col_reg}<16'b1011100100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011100100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100101000000) && ({row_reg, col_reg}<16'b1011100101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011100101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011100101010000) && ({row_reg, col_reg}<16'b1011101001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011101001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101001010111) && ({row_reg, col_reg}<16'b1011101001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011101001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011101001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101001101000) && ({row_reg, col_reg}<16'b1011101010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011101010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101010111011) && ({row_reg, col_reg}<16'b1011101011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011101011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011101011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101011001100) && ({row_reg, col_reg}<16'b1011101100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011101100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101100011011) && ({row_reg, col_reg}<16'b1011101100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011101100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101100101011) && ({row_reg, col_reg}<16'b1011101101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011101101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011101101111101) && ({row_reg, col_reg}<16'b1011101110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011101110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1011101110001101) && ({row_reg, col_reg}<16'b1011110000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011110000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110000011010) && ({row_reg, col_reg}<16'b1011110000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011110000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011110000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110000101011) && ({row_reg, col_reg}<16'b1011110001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011110001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110001111110) && ({row_reg, col_reg}<16'b1011110010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011110010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011110010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110010001111) && ({row_reg, col_reg}<16'b1011110011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011110011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110011011110) && ({row_reg, col_reg}<16'b1011110011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011110011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110011101110) && ({row_reg, col_reg}<16'b1011110100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011110100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110101000000) && ({row_reg, col_reg}<16'b1011110101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011110101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011110101010000) && ({row_reg, col_reg}<16'b1011111001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011111001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111001010111) && ({row_reg, col_reg}<16'b1011111001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011111001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1011111001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111001101000) && ({row_reg, col_reg}<16'b1011111010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011111010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111010111011) && ({row_reg, col_reg}<16'b1011111011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011111011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1011111011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111011001100) && ({row_reg, col_reg}<16'b1011111100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011111100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111100011011) && ({row_reg, col_reg}<16'b1011111100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011111100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111100101011) && ({row_reg, col_reg}<16'b1011111101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1011111101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1011111101111101) && ({row_reg, col_reg}<16'b1011111110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1011111110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1011111110001101) && ({row_reg, col_reg}<16'b1100000000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100000000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000000011010) && ({row_reg, col_reg}<16'b1100000000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100000000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1100000000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000000101011) && ({row_reg, col_reg}<16'b1100000001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100000001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000001111110) && ({row_reg, col_reg}<16'b1100000010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100000010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1100000010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000010001111) && ({row_reg, col_reg}<16'b1100000011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100000011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000011011110) && ({row_reg, col_reg}<16'b1100000011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100000011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000011101110) && ({row_reg, col_reg}<16'b1100000100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100000100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000101000000) && ({row_reg, col_reg}<16'b1100000101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100000101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100000101010000) && ({row_reg, col_reg}<16'b1100001001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100001001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001001010111) && ({row_reg, col_reg}<16'b1100001001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100001001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1100001001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001001101000) && ({row_reg, col_reg}<16'b1100001010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100001010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001010111011) && ({row_reg, col_reg}<16'b1100001011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100001011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1100001011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001011001100) && ({row_reg, col_reg}<16'b1100001100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100001100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001100011011) && ({row_reg, col_reg}<16'b1100001100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100001100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001100101011) && ({row_reg, col_reg}<16'b1100001101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100001101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100001101111101) && ({row_reg, col_reg}<16'b1100001110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100001110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1100001110001101) && ({row_reg, col_reg}<16'b1100010000011001)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100010000011001)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010000011010) && ({row_reg, col_reg}<16'b1100010000101001)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100010000101001)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1100010000101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010000101011) && ({row_reg, col_reg}<16'b1100010001111101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100010001111101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010001111110) && ({row_reg, col_reg}<16'b1100010010001101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100010010001101)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1100010010001110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010010001111) && ({row_reg, col_reg}<16'b1100010011011101)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100010011011101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010011011110) && ({row_reg, col_reg}<16'b1100010011101101)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100010011101101)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010011101110) && ({row_reg, col_reg}<16'b1100010100111111)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100010100111111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010101000000) && ({row_reg, col_reg}<16'b1100010101001111)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100010101001111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100010101010000) && ({row_reg, col_reg}<16'b1100011001010110)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100011001010110)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011001010111) && ({row_reg, col_reg}<16'b1100011001100110)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100011001100110)) color_data = 12'b101110010101;
		if(({row_reg, col_reg}==16'b1100011001100111)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011001101000) && ({row_reg, col_reg}<16'b1100011010111010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100011010111010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011010111011) && ({row_reg, col_reg}<16'b1100011011001010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100011011001010)) color_data = 12'b101110100111;
		if(({row_reg, col_reg}==16'b1100011011001011)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011011001100) && ({row_reg, col_reg}<16'b1100011100011010)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100011100011010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011100011011) && ({row_reg, col_reg}<16'b1100011100101010)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100011100101010)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011100101011) && ({row_reg, col_reg}<16'b1100011101111100)) color_data = 12'b000011110000;
		if(({row_reg, col_reg}==16'b1100011101111100)) color_data = 12'b000000000000;
		if(({row_reg, col_reg}>=16'b1100011101111101) && ({row_reg, col_reg}<16'b1100011110001100)) color_data = 12'b101101110011;
		if(({row_reg, col_reg}==16'b1100011110001100)) color_data = 12'b000000000000;

		if(({row_reg, col_reg}>=16'b1100011110001101) && ({row_reg, col_reg}<16'b1100100000000000)) color_data = 12'b000011110000;

		if(({row_reg, col_reg}>=16'b1100100000000000) && ({row_reg, col_reg}<16'b1100110000000000)) color_data = 12'b000000000000;




		if(({row_reg, col_reg}>=16'b1100110000000000) && ({row_reg, col_reg}<=16'b1101101110011111)) color_data = 12'b000011110000;
	end
endmodule